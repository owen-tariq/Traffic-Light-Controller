library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity My7SegmentDisplay is
port (
        bcd : in std_logic_vector(3 downto 0);  --input
        a, b, c, d, e, f, g : out std_logic;
		  a1, b1, c1, d1, e1, f1, g1 : out std_logic

    );
end My7SegmentDisplay;
--'a' corresponds to MSB of segment7 and g corresponds to LSB of segment7.
architecture Behavioral of My7SegmentDisplay is

begin
process (bcd)
BEGIN
case  bcd is
when "0000" => -- '0'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '0';
		f1 <= '0';
		g1 <= '1';
when "0001"=> -- '1'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '1';
		b1 <= '0';
		c1 <= '0';
		d1 <= '1';
		e1 <= '1';
		f1 <= '1';
		g1 <= '1';
when "0010"=> -- '2'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '1';
		d1 <= '0';
		e1 <= '0';
		f1 <= '1';
		g1 <= '0';
when "0011"=> -- '3'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '1';
		f1 <= '1';
		g1 <= '0';
when "0100"=> -- '4' 
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '1';
		b1 <= '0';
		c1 <= '0';
		d1 <= '1';
		e1 <= '1';
		f1 <= '0';
		g1 <= '0';
when "0101"=> -- '5'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '1';
		c1 <= '0';
		d1 <= '0';
		e1 <= '1';
		f1 <= '0';
		g1 <= '0';
when "0110"=> -- '6'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '1';
		c1 <= '0';
		d1 <= '0';
		e1 <= '0';
		f1 <= '0';
		g1 <= '0';
when "0111"=> -- '7'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '1';
		e1 <= '1';
		f1 <= '1';
		g1 <= '1';
when "1000"=> -- '8'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '0';
		f1 <= '0';
		g1 <= '0';
when "1001"=> -- '9'
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '1';
		f1 <= '0';
		g1 <= '0';
when "1010"=> --'10'
		a <= '1';
		b <= '0';
		c <= '0';
		d <= '1';
		e <= '1';
		f <= '1';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '0';
		f1 <= '0';
		g1 <= '1';
when "1011"=> --'11'
		a <= '1';
		b <= '0';
		c <= '0';
		d <= '1';
		e <= '1';
		f <= '1';
		g <= '1';
		a1 <= '1';
		b1 <= '0';
		c1 <= '0';
		d1 <= '1';
		e1 <= '1';
		f1 <= '1';
		g1 <= '1';
when "1100"=> --'12'
		a <= '1';
		b <= '0';
		c <= '0';
		d <= '1';
		e <= '1';
		f <= '1';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '1';
		d1 <= '0';
		e1 <= '0';
		f1 <= '1';
		g1 <= '0';
when "1101"=> --'13'
		a <= '1';
		b <= '0';
		c <= '0';
		d <= '1';
		e <= '1';
		f <= '1';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '1';
		f1 <= '1';
		g1 <= '0';

when others =>
		a <= '0';
		b <= '0';
		c <= '0';
		d <= '0';
		e <= '0';
		f <= '0';
		g <= '1';
		a1 <= '0';
		b1 <= '0';
		c1 <= '0';
		d1 <= '0';
		e1 <= '0';
		f1 <= '0';
		g1 <= '1';

end case;

end process;

end Behavioral;
